Circuito T2
Vs 1 GND SIN(0 1 1000 0 0 0)
R1 1 2 1.04001336091k
R2 2 5 2.04372276851k
R3 3 2 3.11359737601k
R4 5 GND 4.17085404861k
R5 5 6 3.02859283303k
R6 GND T 2.070545767k
R7 7 8 1.01835949725k
C 6 8 1.00460501759u 
GIb 6 3 (2,5) 7.19043597753m
Vctrl T 7 0V
H1Vd 5 8 Vctrl 8.06397385506k
.ic v(6)=8.765404 v(8)=-1.77636e-15
.end


.control
*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0


echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-5 20e-3

hardcopy trans4.eps v(6) v(1)
echo trans_FIG


quit
.endc

