*
* NGSPICE simulation script
*
*

* forces current values to be saved
.options savecurrents



*Independent Voltage source as transformer
Vs 1 2 SIN(0 21.3386 50 0 0 0)

*envelope detector
D1 1 3 DEF
D2 2 3 DEF
D3 GND 1 DEF
D4 GND 2 DEF
R1 3 GND 150k
C1 3 GND 100u



*voltage regulator
R2 3 4 5k
D5 4 GND D18

.model DEF D
.model D18 D (n=18)
.op
.end

.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0


echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-5 0.6 0.5

***Average***
meas tran yavg AVG v(4) from=500m to=600m

*** max and min vO***
meas tran ymax MAX v(4) from=500m to=600m
meas tran ymin MIN v(4) from=500m to=600m

let vripple = ymax - ymin

print yavg ymax ymin vripple


hardcopy v3.eps v(3)
hardcopy v4.eps  v(4) 
hardcopy v4-12.eps  v(4)-12
echo v3_FIG


quit
.endc
