Circuito T2
.options savecurrents

.INCLUDE ngspice_t23.txt

.ic v(6)=8.765404 v(8)=-1.77636e-15
.op
.end


.control

*makes plots in color
set hcopypscolor=0
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=violet
set color5=rgb:3/8/0
set color6=rgb:4/0/0

echo "********************************************"
echo  "Transient analysis"
echo "********************************************"
tran 1e-5 20e-3

hardcopy trans.eps v(6)
echo trans_FIG


quit
.endc

