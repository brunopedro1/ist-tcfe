Circuito T2
Vs 1 GND 5.20102702949
R1 1 2 1.04001336091k
R2 2 3 2.04372276851k
R3 2 5 3.11359737601k
R4 5 GND 4.17085404861k
R5 5 6 3.02859283303k
R6 GND T 2.070545767k
R7 7 8 1.01835949725k
C 6 8 1.00460501759u 
GIb 6 3 (2,5) 7.19043597753m
Vctrl T 7 0V
H1Vd 5 8 Vctrl 8.06397385506k
.end

.control


op



echo "********************************************"
echo  "Operating point"
echo "********************************************"


echo  "op2_TAB"
print all
echo  "op2_END"




quit
.endc



